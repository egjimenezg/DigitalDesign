----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:52:30 09/06/2014 
-- Module Name:    SIPO - Behavioral 
-- Author:         Gamaliel Jiménez
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SIPO is
    Port ( clock : in  STD_LOGIC);
end SIPO;

architecture Behavioral of SIPO is
begin

end Behavioral;

